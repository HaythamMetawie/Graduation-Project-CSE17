`timescale 1ns / 1ps
`timescale 1ns / 1ps
// This module will be used in weigts generator.
//Generate addresses to get random floating points from randmem.

module random_addresses(output addresses, input wire clk, input wire reset, input wire enable);
	parameter element_width = 32;
	parameter no_of_rand_elements = 16;
	wire [8*no_of_rand_elements - 1:0] addresses; //addresses of random numbers generated by lfsr
	wire up_down = 1; //for lfsr
	wire over_flow; //lfsr overflow output
	genvar i;
	generate
	for(i = 0; i < no_of_rand_elements; i = i +1)
		begin: generate_label
			lfsr my_lfsr(.clk(clk), .resert(reset), .enable(enable), .up_down(up_down), .count(addresses[8*i:8*i + 7]), .overflows(over_flow)); //need to be unique every inst.
		end
	endgenerate		


endmodule
