`timescale 1ns / 1ps
module input_hidden_mem(input wire clk, input wire write_enable, output outData, output reg finish); 

//reg 

endmodule