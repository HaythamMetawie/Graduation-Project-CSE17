`timescale 1ns / 1ps
// This module will be used in weigts generator.

module random_addresses(output addresses, output finish, input wire clk, input wire reset, input wire enable, input read_randMem);
	parameter element_width = 32;
	parameter no_of_rand_elements = 16;
	reg [element_width - 1:0] weigths [0: no_of_rand_elements -1]; //16 random weigths
	reg [7:0] addresses [0: no_of_rand_elements - 1]; //addresses of random numbers generated by lfsr
	wire read_randMem;
	reg finish;
	wire up_down = 1; //for lfsr
	wire over_flow; //lfsr overflow output
	genvar i;
	generate
	for(i = 0; i < no_of_rand_elements; i = i +1)
		begin: generate_label
			lfsr my_lfsr(.clk(clk), .resert(reset), .enable(enable), .up_down(up_down), .count(addresses[j]), .overflows(over_flow)); //need to be unique every inst.
		end
	endgenerate
	
	//random_fp_mem inst(.out_element(weights), .finish(finish), .clk(clk), .addresses(addresses), .readMem(read_randMem));
		


endmodule
